






module control(
clk,



);
input clk;




endmodule