






module control(



)





endmodule