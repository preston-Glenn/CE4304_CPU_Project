






module control(
clk,



)





endmodule