




module Multi_Cycle_Computer(
         clock,
	 reset,
	 program_out
  ) ;
  `include "params.v"

  input clock ;
  input reset ;
  output [DATA_BUS_WIDTH-1:0] program_out ;

  supply1 VDD;













  endmodule